//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2024-04-26
// File Name     : ConvertAB_n4k32_1.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module ConvertAB_n4k32_1(
    input  wire          clk_i,
    input  wire          rst_ni,
    input  wire          i_dvld,
    input  wire          i_rvld,
    input  wire [2559:0] i_n,
    input  wire  [127:0] i_a,
    output wire  [127:0] o_z,
    output wire          o_dvld);

wire     [63:0] x;
wire     [63:0] xd;
wire    [127:0] xp;
wire     [63:0] y;
wire     [63:0] yd;
wire    [127:0] yp;
wire            vrl;
wire            vy;

// ------------------------------------------------------------------------------
// Do ConvertAB(left leaf) instance
// ------------------------------------------------------------------------------
ConvertAB_n2k32_0
  u0_ConvertAB_n2k32_0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[0+:320]),
    .i_a    (i_a[0+:64]),
    .o_z    (x[0+:64]));



// ------------------------------------------------------------------------------
// Connect left leaf data to Expand'input
// ------------------------------------------------------------------------------
assign xd[ 0+:64] = x[ 0+:64];


// ------------------------------------------------------------------------------
// Do a Expand(left leaf) instance
// ------------------------------------------------------------------------------
Expand1_n2o4k32
  u1_Expand1_n2o4k32
   (.i_x  (xd[0+:64]),
    .o_xp (xp[0+:128]));



// ------------------------------------------------------------------------------
// Do ConvertAB(right leaf) instance
// ------------------------------------------------------------------------------
ConvertAB_n2k32_1
  u2_ConvertAB_n2k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[320+:320]),
    .i_a    (i_a[64+:64]),
    .o_z    (y[0+:64]),
    .o_dvld (vrl));



// ------------------------------------------------------------------------------
// Connect right leaf valid to right leaf output
// ------------------------------------------------------------------------------
assign vy = vrl;


// ------------------------------------------------------------------------------
// Connect right leaf data to Expand'input
// ------------------------------------------------------------------------------
assign yd[ 0+:64] = y[ 0+:64];


// ------------------------------------------------------------------------------
// Do a Expand(right leaf) instance
// ------------------------------------------------------------------------------
Expand2_n2o4k32
  u3_Expand2_n2o4k32
   (.i_x  (yd[0+:64]),
    .o_xp (yp[0+:128]));



// ------------------------------------------------------------------------------
// Do a KSA instance
// ------------------------------------------------------------------------------
SecKSA_n4k32_1
  u4_SecKSA_n4k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (vy),
    .i_rvld (i_rvld),
    .i_n    (i_n[640+:1920]),
    .i_x    (xp[0+:128]),
    .i_y    (yp[0+:128]),
    .o_z    (o_z[0+:128]),
    .o_dvld (o_dvld));


endmodule
