//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2023-10-08
// File Name     : SecAnd_PINI1_n2k1_1.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecAnd_PINI1_n2k1_1(
    input  wire       clk_i,
    input  wire       rst_ni,
    input  wire       i_dvld,
    input  wire       i_rvld,
    input  wire [0:0] i_n,
    input  wire [1:0] i_x,
    input  wire [1:0] i_y,
    output wire [1:0] o_c,
    output wire       o_dvld);

(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire  vldd1;// synopsys keep_signal_name "vldd1" 
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xd_0;// synopsys keep_signal_name "xd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xd_1;// synopsys keep_signal_name "xd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yd_0;// synopsys keep_signal_name "yd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yd_1;// synopsys keep_signal_name "yd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_0;// synopsys keep_signal_name "r_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_1;// synopsys keep_signal_name "r_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_0;// synopsys keep_signal_name "yxn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_1;// synopsys keep_signal_name "yxn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_0;// synopsys keep_signal_name "v_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_1;// synopsys keep_signal_name "v_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire vldd2;
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_0;// synopsys keep_signal_name "xdn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_1;// synopsys keep_signal_name "xdn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_0;// synopsys keep_signal_name "xar_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_1;// synopsys keep_signal_name "xar_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_0;// synopsys keep_signal_name "u_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_1;// synopsys keep_signal_name "u_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xay_0;// synopsys keep_signal_name "xay_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xay_1;// synopsys keep_signal_name "xay_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] k_0;// synopsys keep_signal_name "k_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] k_1;// synopsys keep_signal_name "k_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_0;// synopsys keep_signal_name "xav_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_1;// synopsys keep_signal_name "xav_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_0;// synopsys keep_signal_name "t_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_1;// synopsys keep_signal_name "t_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_0;// synopsys keep_signal_name "z_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_1;// synopsys keep_signal_name "z_1"

// delay i_dvld
lix_reg
  #(.W (1))
  u0_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (i_dvld),
    .o_z    (vldd1));



// delay i_x[0+:1]
lix_reg
  #(.W (1))
  u1_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[0+:1]),
    .o_z    (xd_0));



// delay i_x[1+:1]
lix_reg
  #(.W (1))
  u2_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[1+:1]),
    .o_z    (xd_1));



// delay i_y[0+:1]
lix_reg
  #(.W (1))
  u3_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[0+:1]),
    .o_z    (yd_0));



// delay i_y[1+:1]
lix_reg
  #(.W (1))
  u4_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[1+:1]),
    .o_z    (yd_1));



// delay i_n0
lix_reg
  #(.W (1))
  u5_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:1]),
    .o_z    (r_0));



// delay i_n0
lix_reg
  #(.W (1))
  u6_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:1]),
    .o_z    (r_1));



// i_y[0+:1] ^ i_n[0+:1]
lix_xor
  #(.W (1))
  u7_lix_xor
   (.i_x (i_y[1+:1]),
    .i_y (i_n[0+:1]),
    .o_z (yxn_0));



// i_y[1+:1] ^ i_n[0+:1]
lix_xor
  #(.W (1))
  u8_lix_xor
   (.i_x (i_y[0+:1]),
    .i_y (i_n[0+:1]),
    .o_z (yxn_1));



// delay yxn_0
lix_reg
  #(.W (1))
  u9_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_0),
    .o_z    (v_0));



// delay yxn_1
lix_reg
  #(.W (1))
  u10_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_1),
    .o_z    (v_1));



// delay vldd1
lix_reg
  #(.W (1))
  u11_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (vldd1),
    .o_z    (vldd2));



// not  xd_0
lix_not
  #(.W (1))
  u12_lix_not
   (.i_x (xd_0),
    .o_z (xdn_0));



// not  xd_1
lix_not
  #(.W (1))
  u13_lix_not
   (.i_x (xd_1),
    .o_z (xdn_1));



// ~xd_0 & r_0
lix_and
  #(.W (1))
  u14_lix_and
   (.i_x (xdn_0),
    .i_y (r_0),
    .o_z (xar_0));



// ~xd_1 & r_1
lix_and
  #(.W (1))
  u15_lix_and
   (.i_x (xdn_1),
    .i_y (r_1),
    .o_z (xar_1));



// delay ~xd_0 & r_0
lix_reg
  #(.W (1))
  u16_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_0),
    .o_z    (u_0));



// delay ~xd_1 & r_1
lix_reg
  #(.W (1))
  u17_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_1),
    .o_z    (u_1));



// xd_0 & yd_0
lix_and
  #(.W (1))
  u18_lix_and
   (.i_x (xd_0),
    .i_y (yd_0),
    .o_z (xay_0));



// xd_1 & yd_1
lix_and
  #(.W (1))
  u19_lix_and
   (.i_x (xd_1),
    .i_y (yd_1),
    .o_z (xay_1));



// delay xd_0 & yd_0
lix_reg
  #(.W (1))
  u20_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_0),
    .o_z    (k_0));



// delay xd_1 & yd_1
lix_reg
  #(.W (1))
  u21_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_1),
    .o_z    (k_1));



// xd_0 & v_0
lix_and
  #(.W (1))
  u22_lix_and
   (.i_x (xd_0),
    .i_y (v_0),
    .o_z (xav_0));



// xd_1 & v_1
lix_and
  #(.W (1))
  u23_lix_and
   (.i_x (xd_1),
    .i_y (v_1),
    .o_z (xav_1));



// delay xd_0 & v_0
lix_reg
  #(.W (1))
  u24_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_0),
    .o_z    (t_0));



// delay xd_1 & v_1
lix_reg
  #(.W (1))
  u25_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_1),
    .o_z    (t_1));



// u_0 ^ t_0
lix_xor
  #(.W (1))
  u26_lix_xor
   (.i_x (u_0),
    .i_y (t_0),
    .o_z (z_0));



// u_1 ^ t_1
lix_xor
  #(.W (1))
  u27_lix_xor
   (.i_x (u_1),
    .i_y (t_1),
    .o_z (z_1));



// k_0 ^ z_0
lix_xor
  #(.W (1))
  u28_lix_xor
   (.i_x (k_0),
    .i_y (z_0),
    .o_z (o_c[0+:1]));



// k_1 ^ z_1
lix_xor
  #(.W (1))
  u29_lix_xor
   (.i_x (k_1),
    .i_y (z_1),
    .o_z (o_c[1+:1]));



assign o_dvld = vldd2;

endmodule
