//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2023-10-08
// File Name     : SecAnd_PINI1_n5k32_0.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecAnd_PINI1_n5k32_0(
    input  wire         clk_i,
    input  wire         rst_ni,
    input  wire         i_dvld,
    input  wire         i_rvld,
    input  wire [319:0] i_n,
    input  wire [159:0] i_x,
    input  wire [159:0] i_y,
    output wire [159:0] o_c);

(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire  vldd1;// synopsys keep_signal_name "vldd1" 
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_0;// synopsys keep_signal_name "xd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_1;// synopsys keep_signal_name "xd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_2;// synopsys keep_signal_name "xd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_3;// synopsys keep_signal_name "xd_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_4;// synopsys keep_signal_name "xd_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_0;// synopsys keep_signal_name "yd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_1;// synopsys keep_signal_name "yd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_2;// synopsys keep_signal_name "yd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_3;// synopsys keep_signal_name "yd_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_4;// synopsys keep_signal_name "yd_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_0;// synopsys keep_signal_name "r_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_1;// synopsys keep_signal_name "r_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_2;// synopsys keep_signal_name "r_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_3;// synopsys keep_signal_name "r_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_4;// synopsys keep_signal_name "r_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_5;// synopsys keep_signal_name "r_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_6;// synopsys keep_signal_name "r_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_7;// synopsys keep_signal_name "r_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_8;// synopsys keep_signal_name "r_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_9;// synopsys keep_signal_name "r_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_10;// synopsys keep_signal_name "r_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_11;// synopsys keep_signal_name "r_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_12;// synopsys keep_signal_name "r_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_13;// synopsys keep_signal_name "r_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_14;// synopsys keep_signal_name "r_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_15;// synopsys keep_signal_name "r_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_16;// synopsys keep_signal_name "r_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_17;// synopsys keep_signal_name "r_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_18;// synopsys keep_signal_name "r_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_19;// synopsys keep_signal_name "r_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_0;// synopsys keep_signal_name "yxn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_1;// synopsys keep_signal_name "yxn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_2;// synopsys keep_signal_name "yxn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_3;// synopsys keep_signal_name "yxn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_4;// synopsys keep_signal_name "yxn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_5;// synopsys keep_signal_name "yxn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_6;// synopsys keep_signal_name "yxn_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_7;// synopsys keep_signal_name "yxn_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_8;// synopsys keep_signal_name "yxn_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_9;// synopsys keep_signal_name "yxn_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_10;// synopsys keep_signal_name "yxn_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_11;// synopsys keep_signal_name "yxn_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_12;// synopsys keep_signal_name "yxn_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_13;// synopsys keep_signal_name "yxn_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_14;// synopsys keep_signal_name "yxn_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_15;// synopsys keep_signal_name "yxn_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_16;// synopsys keep_signal_name "yxn_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_17;// synopsys keep_signal_name "yxn_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_18;// synopsys keep_signal_name "yxn_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_19;// synopsys keep_signal_name "yxn_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_0;// synopsys keep_signal_name "v_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_1;// synopsys keep_signal_name "v_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_2;// synopsys keep_signal_name "v_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_3;// synopsys keep_signal_name "v_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_4;// synopsys keep_signal_name "v_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_5;// synopsys keep_signal_name "v_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_6;// synopsys keep_signal_name "v_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_7;// synopsys keep_signal_name "v_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_8;// synopsys keep_signal_name "v_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_9;// synopsys keep_signal_name "v_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_10;// synopsys keep_signal_name "v_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_11;// synopsys keep_signal_name "v_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_12;// synopsys keep_signal_name "v_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_13;// synopsys keep_signal_name "v_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_14;// synopsys keep_signal_name "v_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_15;// synopsys keep_signal_name "v_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_16;// synopsys keep_signal_name "v_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_17;// synopsys keep_signal_name "v_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_18;// synopsys keep_signal_name "v_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_19;// synopsys keep_signal_name "v_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_0;// synopsys keep_signal_name "xdn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_1;// synopsys keep_signal_name "xdn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_2;// synopsys keep_signal_name "xdn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_3;// synopsys keep_signal_name "xdn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_4;// synopsys keep_signal_name "xdn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_5;// synopsys keep_signal_name "xdn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_6;// synopsys keep_signal_name "xdn_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_7;// synopsys keep_signal_name "xdn_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_8;// synopsys keep_signal_name "xdn_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_9;// synopsys keep_signal_name "xdn_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_10;// synopsys keep_signal_name "xdn_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_11;// synopsys keep_signal_name "xdn_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_12;// synopsys keep_signal_name "xdn_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_13;// synopsys keep_signal_name "xdn_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_14;// synopsys keep_signal_name "xdn_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_15;// synopsys keep_signal_name "xdn_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_16;// synopsys keep_signal_name "xdn_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_17;// synopsys keep_signal_name "xdn_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_18;// synopsys keep_signal_name "xdn_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_19;// synopsys keep_signal_name "xdn_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_0;// synopsys keep_signal_name "xar_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_1;// synopsys keep_signal_name "xar_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_2;// synopsys keep_signal_name "xar_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_3;// synopsys keep_signal_name "xar_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_4;// synopsys keep_signal_name "xar_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_5;// synopsys keep_signal_name "xar_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_6;// synopsys keep_signal_name "xar_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_7;// synopsys keep_signal_name "xar_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_8;// synopsys keep_signal_name "xar_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_9;// synopsys keep_signal_name "xar_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_10;// synopsys keep_signal_name "xar_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_11;// synopsys keep_signal_name "xar_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_12;// synopsys keep_signal_name "xar_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_13;// synopsys keep_signal_name "xar_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_14;// synopsys keep_signal_name "xar_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_15;// synopsys keep_signal_name "xar_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_16;// synopsys keep_signal_name "xar_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_17;// synopsys keep_signal_name "xar_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_18;// synopsys keep_signal_name "xar_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_19;// synopsys keep_signal_name "xar_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_0;// synopsys keep_signal_name "u_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_1;// synopsys keep_signal_name "u_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_2;// synopsys keep_signal_name "u_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_3;// synopsys keep_signal_name "u_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_4;// synopsys keep_signal_name "u_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_5;// synopsys keep_signal_name "u_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_6;// synopsys keep_signal_name "u_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_7;// synopsys keep_signal_name "u_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_8;// synopsys keep_signal_name "u_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_9;// synopsys keep_signal_name "u_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_10;// synopsys keep_signal_name "u_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_11;// synopsys keep_signal_name "u_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_12;// synopsys keep_signal_name "u_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_13;// synopsys keep_signal_name "u_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_14;// synopsys keep_signal_name "u_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_15;// synopsys keep_signal_name "u_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_16;// synopsys keep_signal_name "u_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_17;// synopsys keep_signal_name "u_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_18;// synopsys keep_signal_name "u_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_19;// synopsys keep_signal_name "u_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_0;// synopsys keep_signal_name "xay_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_1;// synopsys keep_signal_name "xay_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_2;// synopsys keep_signal_name "xay_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_3;// synopsys keep_signal_name "xay_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_4;// synopsys keep_signal_name "xay_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_0;// synopsys keep_signal_name "k_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_1;// synopsys keep_signal_name "k_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_2;// synopsys keep_signal_name "k_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_3;// synopsys keep_signal_name "k_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_4;// synopsys keep_signal_name "k_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_0;// synopsys keep_signal_name "xav_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_1;// synopsys keep_signal_name "xav_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_2;// synopsys keep_signal_name "xav_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_3;// synopsys keep_signal_name "xav_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_4;// synopsys keep_signal_name "xav_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_5;// synopsys keep_signal_name "xav_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_6;// synopsys keep_signal_name "xav_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_7;// synopsys keep_signal_name "xav_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_8;// synopsys keep_signal_name "xav_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_9;// synopsys keep_signal_name "xav_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_10;// synopsys keep_signal_name "xav_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_11;// synopsys keep_signal_name "xav_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_12;// synopsys keep_signal_name "xav_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_13;// synopsys keep_signal_name "xav_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_14;// synopsys keep_signal_name "xav_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_15;// synopsys keep_signal_name "xav_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_16;// synopsys keep_signal_name "xav_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_17;// synopsys keep_signal_name "xav_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_18;// synopsys keep_signal_name "xav_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_19;// synopsys keep_signal_name "xav_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_0;// synopsys keep_signal_name "t_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_1;// synopsys keep_signal_name "t_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_2;// synopsys keep_signal_name "t_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_3;// synopsys keep_signal_name "t_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_4;// synopsys keep_signal_name "t_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_5;// synopsys keep_signal_name "t_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_6;// synopsys keep_signal_name "t_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_7;// synopsys keep_signal_name "t_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_8;// synopsys keep_signal_name "t_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_9;// synopsys keep_signal_name "t_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_10;// synopsys keep_signal_name "t_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_11;// synopsys keep_signal_name "t_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_12;// synopsys keep_signal_name "t_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_13;// synopsys keep_signal_name "t_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_14;// synopsys keep_signal_name "t_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_15;// synopsys keep_signal_name "t_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_16;// synopsys keep_signal_name "t_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_17;// synopsys keep_signal_name "t_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_18;// synopsys keep_signal_name "t_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_19;// synopsys keep_signal_name "t_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_0;// synopsys keep_signal_name "z_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_1;// synopsys keep_signal_name "z_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_2;// synopsys keep_signal_name "z_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_3;// synopsys keep_signal_name "z_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_4;// synopsys keep_signal_name "z_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_5;// synopsys keep_signal_name "z_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_6;// synopsys keep_signal_name "z_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_7;// synopsys keep_signal_name "z_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_8;// synopsys keep_signal_name "z_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_9;// synopsys keep_signal_name "z_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_10;// synopsys keep_signal_name "z_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_11;// synopsys keep_signal_name "z_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_12;// synopsys keep_signal_name "z_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_13;// synopsys keep_signal_name "z_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_14;// synopsys keep_signal_name "z_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_15;// synopsys keep_signal_name "z_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_16;// synopsys keep_signal_name "z_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_17;// synopsys keep_signal_name "z_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_18;// synopsys keep_signal_name "z_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_19;// synopsys keep_signal_name "z_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_0;// synopsys keep_signal_name "zxz_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_1;// synopsys keep_signal_name "zxz_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_2;// synopsys keep_signal_name "zxz_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_3;// synopsys keep_signal_name "zxz_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_4;// synopsys keep_signal_name "zxz_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_5;// synopsys keep_signal_name "zxz_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_6;// synopsys keep_signal_name "zxz_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_7;// synopsys keep_signal_name "zxz_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_8;// synopsys keep_signal_name "zxz_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_9;// synopsys keep_signal_name "zxz_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_10;// synopsys keep_signal_name "zxz_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_11;// synopsys keep_signal_name "zxz_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_12;// synopsys keep_signal_name "zxz_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_13;// synopsys keep_signal_name "zxz_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_14;// synopsys keep_signal_name "zxz_14"

// delay i_dvld
lix_reg
  #(.W (1))
  u0_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (i_dvld),
    .o_z    (vldd1));



// delay i_x[0+:32]
lix_reg
  #(.W (32))
  u1_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[0+:32]),
    .o_z    (xd_0));



// delay i_x[32+:32]
lix_reg
  #(.W (32))
  u2_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[32+:32]),
    .o_z    (xd_1));



// delay i_x[64+:32]
lix_reg
  #(.W (32))
  u3_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[64+:32]),
    .o_z    (xd_2));



// delay i_x[96+:32]
lix_reg
  #(.W (32))
  u4_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[96+:32]),
    .o_z    (xd_3));



// delay i_x[128+:32]
lix_reg
  #(.W (32))
  u5_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[128+:32]),
    .o_z    (xd_4));



// delay i_y[0+:32]
lix_reg
  #(.W (32))
  u6_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[0+:32]),
    .o_z    (yd_0));



// delay i_y[32+:32]
lix_reg
  #(.W (32))
  u7_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[32+:32]),
    .o_z    (yd_1));



// delay i_y[64+:32]
lix_reg
  #(.W (32))
  u8_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[64+:32]),
    .o_z    (yd_2));



// delay i_y[96+:32]
lix_reg
  #(.W (32))
  u9_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[96+:32]),
    .o_z    (yd_3));



// delay i_y[128+:32]
lix_reg
  #(.W (32))
  u10_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[128+:32]),
    .o_z    (yd_4));



// delay i_n0
lix_reg
  #(.W (32))
  u11_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:32]),
    .o_z    (r_0));



// delay i_n1
lix_reg
  #(.W (32))
  u12_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[32+:32]),
    .o_z    (r_1));



// delay i_n2
lix_reg
  #(.W (32))
  u13_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[64+:32]),
    .o_z    (r_2));



// delay i_n3
lix_reg
  #(.W (32))
  u14_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[96+:32]),
    .o_z    (r_3));



// delay i_n0
lix_reg
  #(.W (32))
  u15_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:32]),
    .o_z    (r_4));



// delay i_n4
lix_reg
  #(.W (32))
  u16_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[128+:32]),
    .o_z    (r_5));



// delay i_n5
lix_reg
  #(.W (32))
  u17_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[160+:32]),
    .o_z    (r_6));



// delay i_n6
lix_reg
  #(.W (32))
  u18_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[192+:32]),
    .o_z    (r_7));



// delay i_n1
lix_reg
  #(.W (32))
  u19_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[32+:32]),
    .o_z    (r_8));



// delay i_n4
lix_reg
  #(.W (32))
  u20_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[128+:32]),
    .o_z    (r_9));



// delay i_n7
lix_reg
  #(.W (32))
  u21_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[224+:32]),
    .o_z    (r_10));



// delay i_n8
lix_reg
  #(.W (32))
  u22_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[256+:32]),
    .o_z    (r_11));



// delay i_n2
lix_reg
  #(.W (32))
  u23_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[64+:32]),
    .o_z    (r_12));



// delay i_n5
lix_reg
  #(.W (32))
  u24_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[160+:32]),
    .o_z    (r_13));



// delay i_n7
lix_reg
  #(.W (32))
  u25_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[224+:32]),
    .o_z    (r_14));



// delay i_n9
lix_reg
  #(.W (32))
  u26_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[288+:32]),
    .o_z    (r_15));



// delay i_n3
lix_reg
  #(.W (32))
  u27_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[96+:32]),
    .o_z    (r_16));



// delay i_n6
lix_reg
  #(.W (32))
  u28_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[192+:32]),
    .o_z    (r_17));



// delay i_n8
lix_reg
  #(.W (32))
  u29_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[256+:32]),
    .o_z    (r_18));



// delay i_n9
lix_reg
  #(.W (32))
  u30_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[288+:32]),
    .o_z    (r_19));



// i_y[0+:32] ^ i_n[0+:32]
lix_xor
  #(.W (32))
  u31_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[0+:32]),
    .o_z (yxn_0));



// i_y[0+:32] ^ i_n[32+:32]
lix_xor
  #(.W (32))
  u32_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[32+:32]),
    .o_z (yxn_1));



// i_y[0+:32] ^ i_n[64+:32]
lix_xor
  #(.W (32))
  u33_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[64+:32]),
    .o_z (yxn_2));



// i_y[0+:32] ^ i_n[96+:32]
lix_xor
  #(.W (32))
  u34_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[96+:32]),
    .o_z (yxn_3));



// i_y[32+:32] ^ i_n[0+:32]
lix_xor
  #(.W (32))
  u35_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[0+:32]),
    .o_z (yxn_4));



// i_y[32+:32] ^ i_n[128+:32]
lix_xor
  #(.W (32))
  u36_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[128+:32]),
    .o_z (yxn_5));



// i_y[32+:32] ^ i_n[160+:32]
lix_xor
  #(.W (32))
  u37_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[160+:32]),
    .o_z (yxn_6));



// i_y[32+:32] ^ i_n[192+:32]
lix_xor
  #(.W (32))
  u38_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[192+:32]),
    .o_z (yxn_7));



// i_y[64+:32] ^ i_n[32+:32]
lix_xor
  #(.W (32))
  u39_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[32+:32]),
    .o_z (yxn_8));



// i_y[64+:32] ^ i_n[128+:32]
lix_xor
  #(.W (32))
  u40_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[128+:32]),
    .o_z (yxn_9));



// i_y[64+:32] ^ i_n[224+:32]
lix_xor
  #(.W (32))
  u41_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[224+:32]),
    .o_z (yxn_10));



// i_y[64+:32] ^ i_n[256+:32]
lix_xor
  #(.W (32))
  u42_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[256+:32]),
    .o_z (yxn_11));



// i_y[96+:32] ^ i_n[64+:32]
lix_xor
  #(.W (32))
  u43_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[64+:32]),
    .o_z (yxn_12));



// i_y[96+:32] ^ i_n[160+:32]
lix_xor
  #(.W (32))
  u44_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[160+:32]),
    .o_z (yxn_13));



// i_y[96+:32] ^ i_n[224+:32]
lix_xor
  #(.W (32))
  u45_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[224+:32]),
    .o_z (yxn_14));



// i_y[96+:32] ^ i_n[288+:32]
lix_xor
  #(.W (32))
  u46_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[288+:32]),
    .o_z (yxn_15));



// i_y[128+:32] ^ i_n[96+:32]
lix_xor
  #(.W (32))
  u47_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[96+:32]),
    .o_z (yxn_16));



// i_y[128+:32] ^ i_n[192+:32]
lix_xor
  #(.W (32))
  u48_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[192+:32]),
    .o_z (yxn_17));



// i_y[128+:32] ^ i_n[256+:32]
lix_xor
  #(.W (32))
  u49_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[256+:32]),
    .o_z (yxn_18));



// i_y[128+:32] ^ i_n[288+:32]
lix_xor
  #(.W (32))
  u50_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[288+:32]),
    .o_z (yxn_19));



// delay yxn_0
lix_reg
  #(.W (32))
  u51_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_0),
    .o_z    (v_0));



// delay yxn_1
lix_reg
  #(.W (32))
  u52_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_1),
    .o_z    (v_1));



// delay yxn_2
lix_reg
  #(.W (32))
  u53_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_2),
    .o_z    (v_2));



// delay yxn_3
lix_reg
  #(.W (32))
  u54_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_3),
    .o_z    (v_3));



// delay yxn_4
lix_reg
  #(.W (32))
  u55_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_4),
    .o_z    (v_4));



// delay yxn_5
lix_reg
  #(.W (32))
  u56_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_5),
    .o_z    (v_5));



// delay yxn_6
lix_reg
  #(.W (32))
  u57_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_6),
    .o_z    (v_6));



// delay yxn_7
lix_reg
  #(.W (32))
  u58_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_7),
    .o_z    (v_7));



// delay yxn_8
lix_reg
  #(.W (32))
  u59_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_8),
    .o_z    (v_8));



// delay yxn_9
lix_reg
  #(.W (32))
  u60_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_9),
    .o_z    (v_9));



// delay yxn_10
lix_reg
  #(.W (32))
  u61_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_10),
    .o_z    (v_10));



// delay yxn_11
lix_reg
  #(.W (32))
  u62_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_11),
    .o_z    (v_11));



// delay yxn_12
lix_reg
  #(.W (32))
  u63_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_12),
    .o_z    (v_12));



// delay yxn_13
lix_reg
  #(.W (32))
  u64_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_13),
    .o_z    (v_13));



// delay yxn_14
lix_reg
  #(.W (32))
  u65_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_14),
    .o_z    (v_14));



// delay yxn_15
lix_reg
  #(.W (32))
  u66_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_15),
    .o_z    (v_15));



// delay yxn_16
lix_reg
  #(.W (32))
  u67_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_16),
    .o_z    (v_16));



// delay yxn_17
lix_reg
  #(.W (32))
  u68_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_17),
    .o_z    (v_17));



// delay yxn_18
lix_reg
  #(.W (32))
  u69_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_18),
    .o_z    (v_18));



// delay yxn_19
lix_reg
  #(.W (32))
  u70_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_19),
    .o_z    (v_19));



// not  xd_0
lix_not
  #(.W (32))
  u71_lix_not
   (.i_x (xd_0),
    .o_z (xdn_0));



// not  xd_1
lix_not
  #(.W (32))
  u72_lix_not
   (.i_x (xd_1),
    .o_z (xdn_1));



// not  xd_2
lix_not
  #(.W (32))
  u73_lix_not
   (.i_x (xd_2),
    .o_z (xdn_2));



// not  xd_3
lix_not
  #(.W (32))
  u74_lix_not
   (.i_x (xd_3),
    .o_z (xdn_3));



// not  xd_4
lix_not
  #(.W (32))
  u75_lix_not
   (.i_x (xd_4),
    .o_z (xdn_4));



// ~xd_0 & r_0
lix_and
  #(.W (32))
  u76_lix_and
   (.i_x (xdn_0),
    .i_y (r_0),
    .o_z (xar_0));



// ~xd_0 & r_1
lix_and
  #(.W (32))
  u77_lix_and
   (.i_x (xdn_0),
    .i_y (r_1),
    .o_z (xar_1));



// ~xd_0 & r_2
lix_and
  #(.W (32))
  u78_lix_and
   (.i_x (xdn_0),
    .i_y (r_2),
    .o_z (xar_2));



// ~xd_0 & r_3
lix_and
  #(.W (32))
  u79_lix_and
   (.i_x (xdn_0),
    .i_y (r_3),
    .o_z (xar_3));



// ~xd_1 & r_4
lix_and
  #(.W (32))
  u80_lix_and
   (.i_x (xdn_1),
    .i_y (r_4),
    .o_z (xar_4));



// ~xd_1 & r_5
lix_and
  #(.W (32))
  u81_lix_and
   (.i_x (xdn_1),
    .i_y (r_5),
    .o_z (xar_5));



// ~xd_1 & r_6
lix_and
  #(.W (32))
  u82_lix_and
   (.i_x (xdn_1),
    .i_y (r_6),
    .o_z (xar_6));



// ~xd_1 & r_7
lix_and
  #(.W (32))
  u83_lix_and
   (.i_x (xdn_1),
    .i_y (r_7),
    .o_z (xar_7));



// ~xd_2 & r_8
lix_and
  #(.W (32))
  u84_lix_and
   (.i_x (xdn_2),
    .i_y (r_8),
    .o_z (xar_8));



// ~xd_2 & r_9
lix_and
  #(.W (32))
  u85_lix_and
   (.i_x (xdn_2),
    .i_y (r_9),
    .o_z (xar_9));



// ~xd_2 & r_10
lix_and
  #(.W (32))
  u86_lix_and
   (.i_x (xdn_2),
    .i_y (r_10),
    .o_z (xar_10));



// ~xd_2 & r_11
lix_and
  #(.W (32))
  u87_lix_and
   (.i_x (xdn_2),
    .i_y (r_11),
    .o_z (xar_11));



// ~xd_3 & r_12
lix_and
  #(.W (32))
  u88_lix_and
   (.i_x (xdn_3),
    .i_y (r_12),
    .o_z (xar_12));



// ~xd_3 & r_13
lix_and
  #(.W (32))
  u89_lix_and
   (.i_x (xdn_3),
    .i_y (r_13),
    .o_z (xar_13));



// ~xd_3 & r_14
lix_and
  #(.W (32))
  u90_lix_and
   (.i_x (xdn_3),
    .i_y (r_14),
    .o_z (xar_14));



// ~xd_3 & r_15
lix_and
  #(.W (32))
  u91_lix_and
   (.i_x (xdn_3),
    .i_y (r_15),
    .o_z (xar_15));



// ~xd_4 & r_16
lix_and
  #(.W (32))
  u92_lix_and
   (.i_x (xdn_4),
    .i_y (r_16),
    .o_z (xar_16));



// ~xd_4 & r_17
lix_and
  #(.W (32))
  u93_lix_and
   (.i_x (xdn_4),
    .i_y (r_17),
    .o_z (xar_17));



// ~xd_4 & r_18
lix_and
  #(.W (32))
  u94_lix_and
   (.i_x (xdn_4),
    .i_y (r_18),
    .o_z (xar_18));



// ~xd_4 & r_19
lix_and
  #(.W (32))
  u95_lix_and
   (.i_x (xdn_4),
    .i_y (r_19),
    .o_z (xar_19));



// delay ~xd_0 & r_0
lix_reg
  #(.W (32))
  u96_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_0),
    .o_z    (u_0));



// delay ~xd_1 & r_1
lix_reg
  #(.W (32))
  u97_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_1),
    .o_z    (u_1));



// delay ~xd_2 & r_2
lix_reg
  #(.W (32))
  u98_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_2),
    .o_z    (u_2));



// delay ~xd_3 & r_3
lix_reg
  #(.W (32))
  u99_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_3),
    .o_z    (u_3));



// delay ~xd_4 & r_4
lix_reg
  #(.W (32))
  u100_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_4),
    .o_z    (u_4));



// delay ~xd_5 & r_5
lix_reg
  #(.W (32))
  u101_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_5),
    .o_z    (u_5));



// delay ~xd_6 & r_6
lix_reg
  #(.W (32))
  u102_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_6),
    .o_z    (u_6));



// delay ~xd_7 & r_7
lix_reg
  #(.W (32))
  u103_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_7),
    .o_z    (u_7));



// delay ~xd_8 & r_8
lix_reg
  #(.W (32))
  u104_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_8),
    .o_z    (u_8));



// delay ~xd_9 & r_9
lix_reg
  #(.W (32))
  u105_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_9),
    .o_z    (u_9));



// delay ~xd_10 & r_10
lix_reg
  #(.W (32))
  u106_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_10),
    .o_z    (u_10));



// delay ~xd_11 & r_11
lix_reg
  #(.W (32))
  u107_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_11),
    .o_z    (u_11));



// delay ~xd_12 & r_12
lix_reg
  #(.W (32))
  u108_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_12),
    .o_z    (u_12));



// delay ~xd_13 & r_13
lix_reg
  #(.W (32))
  u109_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_13),
    .o_z    (u_13));



// delay ~xd_14 & r_14
lix_reg
  #(.W (32))
  u110_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_14),
    .o_z    (u_14));



// delay ~xd_15 & r_15
lix_reg
  #(.W (32))
  u111_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_15),
    .o_z    (u_15));



// delay ~xd_16 & r_16
lix_reg
  #(.W (32))
  u112_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_16),
    .o_z    (u_16));



// delay ~xd_17 & r_17
lix_reg
  #(.W (32))
  u113_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_17),
    .o_z    (u_17));



// delay ~xd_18 & r_18
lix_reg
  #(.W (32))
  u114_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_18),
    .o_z    (u_18));



// delay ~xd_19 & r_19
lix_reg
  #(.W (32))
  u115_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_19),
    .o_z    (u_19));



// xd_0 & yd_0
lix_and
  #(.W (32))
  u116_lix_and
   (.i_x (xd_0),
    .i_y (yd_0),
    .o_z (xay_0));



// xd_1 & yd_1
lix_and
  #(.W (32))
  u117_lix_and
   (.i_x (xd_1),
    .i_y (yd_1),
    .o_z (xay_1));



// xd_2 & yd_2
lix_and
  #(.W (32))
  u118_lix_and
   (.i_x (xd_2),
    .i_y (yd_2),
    .o_z (xay_2));



// xd_3 & yd_3
lix_and
  #(.W (32))
  u119_lix_and
   (.i_x (xd_3),
    .i_y (yd_3),
    .o_z (xay_3));



// xd_4 & yd_4
lix_and
  #(.W (32))
  u120_lix_and
   (.i_x (xd_4),
    .i_y (yd_4),
    .o_z (xay_4));



// delay xd_0 & yd_0
lix_reg
  #(.W (32))
  u121_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_0),
    .o_z    (k_0));



// delay xd_1 & yd_1
lix_reg
  #(.W (32))
  u122_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_1),
    .o_z    (k_1));



// delay xd_2 & yd_2
lix_reg
  #(.W (32))
  u123_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_2),
    .o_z    (k_2));



// delay xd_3 & yd_3
lix_reg
  #(.W (32))
  u124_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_3),
    .o_z    (k_3));



// delay xd_4 & yd_4
lix_reg
  #(.W (32))
  u125_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_4),
    .o_z    (k_4));



// xd_0 & v_0
lix_and
  #(.W (32))
  u126_lix_and
   (.i_x (xd_0),
    .i_y (v_0),
    .o_z (xav_0));



// xd_0 & v_1
lix_and
  #(.W (32))
  u127_lix_and
   (.i_x (xd_0),
    .i_y (v_1),
    .o_z (xav_1));



// xd_0 & v_2
lix_and
  #(.W (32))
  u128_lix_and
   (.i_x (xd_0),
    .i_y (v_2),
    .o_z (xav_2));



// xd_0 & v_3
lix_and
  #(.W (32))
  u129_lix_and
   (.i_x (xd_0),
    .i_y (v_3),
    .o_z (xav_3));



// xd_1 & v_4
lix_and
  #(.W (32))
  u130_lix_and
   (.i_x (xd_1),
    .i_y (v_4),
    .o_z (xav_4));



// xd_1 & v_5
lix_and
  #(.W (32))
  u131_lix_and
   (.i_x (xd_1),
    .i_y (v_5),
    .o_z (xav_5));



// xd_1 & v_6
lix_and
  #(.W (32))
  u132_lix_and
   (.i_x (xd_1),
    .i_y (v_6),
    .o_z (xav_6));



// xd_1 & v_7
lix_and
  #(.W (32))
  u133_lix_and
   (.i_x (xd_1),
    .i_y (v_7),
    .o_z (xav_7));



// xd_2 & v_8
lix_and
  #(.W (32))
  u134_lix_and
   (.i_x (xd_2),
    .i_y (v_8),
    .o_z (xav_8));



// xd_2 & v_9
lix_and
  #(.W (32))
  u135_lix_and
   (.i_x (xd_2),
    .i_y (v_9),
    .o_z (xav_9));



// xd_2 & v_10
lix_and
  #(.W (32))
  u136_lix_and
   (.i_x (xd_2),
    .i_y (v_10),
    .o_z (xav_10));



// xd_2 & v_11
lix_and
  #(.W (32))
  u137_lix_and
   (.i_x (xd_2),
    .i_y (v_11),
    .o_z (xav_11));



// xd_3 & v_12
lix_and
  #(.W (32))
  u138_lix_and
   (.i_x (xd_3),
    .i_y (v_12),
    .o_z (xav_12));



// xd_3 & v_13
lix_and
  #(.W (32))
  u139_lix_and
   (.i_x (xd_3),
    .i_y (v_13),
    .o_z (xav_13));



// xd_3 & v_14
lix_and
  #(.W (32))
  u140_lix_and
   (.i_x (xd_3),
    .i_y (v_14),
    .o_z (xav_14));



// xd_3 & v_15
lix_and
  #(.W (32))
  u141_lix_and
   (.i_x (xd_3),
    .i_y (v_15),
    .o_z (xav_15));



// xd_4 & v_16
lix_and
  #(.W (32))
  u142_lix_and
   (.i_x (xd_4),
    .i_y (v_16),
    .o_z (xav_16));



// xd_4 & v_17
lix_and
  #(.W (32))
  u143_lix_and
   (.i_x (xd_4),
    .i_y (v_17),
    .o_z (xav_17));



// xd_4 & v_18
lix_and
  #(.W (32))
  u144_lix_and
   (.i_x (xd_4),
    .i_y (v_18),
    .o_z (xav_18));



// xd_4 & v_19
lix_and
  #(.W (32))
  u145_lix_and
   (.i_x (xd_4),
    .i_y (v_19),
    .o_z (xav_19));



// delay xd_0 & v_0
lix_reg
  #(.W (32))
  u146_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_0),
    .o_z    (t_0));



// delay xd_1 & v_1
lix_reg
  #(.W (32))
  u147_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_1),
    .o_z    (t_1));



// delay xd_2 & v_2
lix_reg
  #(.W (32))
  u148_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_2),
    .o_z    (t_2));



// delay xd_3 & v_3
lix_reg
  #(.W (32))
  u149_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_3),
    .o_z    (t_3));



// delay xd_4 & v_4
lix_reg
  #(.W (32))
  u150_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_4),
    .o_z    (t_4));



// delay xd_5 & v_5
lix_reg
  #(.W (32))
  u151_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_5),
    .o_z    (t_5));



// delay xd_6 & v_6
lix_reg
  #(.W (32))
  u152_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_6),
    .o_z    (t_6));



// delay xd_7 & v_7
lix_reg
  #(.W (32))
  u153_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_7),
    .o_z    (t_7));



// delay xd_8 & v_8
lix_reg
  #(.W (32))
  u154_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_8),
    .o_z    (t_8));



// delay xd_9 & v_9
lix_reg
  #(.W (32))
  u155_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_9),
    .o_z    (t_9));



// delay xd_10 & v_10
lix_reg
  #(.W (32))
  u156_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_10),
    .o_z    (t_10));



// delay xd_11 & v_11
lix_reg
  #(.W (32))
  u157_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_11),
    .o_z    (t_11));



// delay xd_12 & v_12
lix_reg
  #(.W (32))
  u158_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_12),
    .o_z    (t_12));



// delay xd_13 & v_13
lix_reg
  #(.W (32))
  u159_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_13),
    .o_z    (t_13));



// delay xd_14 & v_14
lix_reg
  #(.W (32))
  u160_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_14),
    .o_z    (t_14));



// delay xd_15 & v_15
lix_reg
  #(.W (32))
  u161_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_15),
    .o_z    (t_15));



// delay xd_16 & v_16
lix_reg
  #(.W (32))
  u162_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_16),
    .o_z    (t_16));



// delay xd_17 & v_17
lix_reg
  #(.W (32))
  u163_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_17),
    .o_z    (t_17));



// delay xd_18 & v_18
lix_reg
  #(.W (32))
  u164_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_18),
    .o_z    (t_18));



// delay xd_19 & v_19
lix_reg
  #(.W (32))
  u165_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_19),
    .o_z    (t_19));



// u_0 ^ t_0
lix_xor
  #(.W (32))
  u166_lix_xor
   (.i_x (u_0),
    .i_y (t_0),
    .o_z (z_0));



// u_1 ^ t_1
lix_xor
  #(.W (32))
  u167_lix_xor
   (.i_x (u_1),
    .i_y (t_1),
    .o_z (z_1));



// u_2 ^ t_2
lix_xor
  #(.W (32))
  u168_lix_xor
   (.i_x (u_2),
    .i_y (t_2),
    .o_z (z_2));



// u_3 ^ t_3
lix_xor
  #(.W (32))
  u169_lix_xor
   (.i_x (u_3),
    .i_y (t_3),
    .o_z (z_3));



// u_4 ^ t_4
lix_xor
  #(.W (32))
  u170_lix_xor
   (.i_x (u_4),
    .i_y (t_4),
    .o_z (z_4));



// u_5 ^ t_5
lix_xor
  #(.W (32))
  u171_lix_xor
   (.i_x (u_5),
    .i_y (t_5),
    .o_z (z_5));



// u_6 ^ t_6
lix_xor
  #(.W (32))
  u172_lix_xor
   (.i_x (u_6),
    .i_y (t_6),
    .o_z (z_6));



// u_7 ^ t_7
lix_xor
  #(.W (32))
  u173_lix_xor
   (.i_x (u_7),
    .i_y (t_7),
    .o_z (z_7));



// u_8 ^ t_8
lix_xor
  #(.W (32))
  u174_lix_xor
   (.i_x (u_8),
    .i_y (t_8),
    .o_z (z_8));



// u_9 ^ t_9
lix_xor
  #(.W (32))
  u175_lix_xor
   (.i_x (u_9),
    .i_y (t_9),
    .o_z (z_9));



// u_10 ^ t_10
lix_xor
  #(.W (32))
  u176_lix_xor
   (.i_x (u_10),
    .i_y (t_10),
    .o_z (z_10));



// u_11 ^ t_11
lix_xor
  #(.W (32))
  u177_lix_xor
   (.i_x (u_11),
    .i_y (t_11),
    .o_z (z_11));



// u_12 ^ t_12
lix_xor
  #(.W (32))
  u178_lix_xor
   (.i_x (u_12),
    .i_y (t_12),
    .o_z (z_12));



// u_13 ^ t_13
lix_xor
  #(.W (32))
  u179_lix_xor
   (.i_x (u_13),
    .i_y (t_13),
    .o_z (z_13));



// u_14 ^ t_14
lix_xor
  #(.W (32))
  u180_lix_xor
   (.i_x (u_14),
    .i_y (t_14),
    .o_z (z_14));



// u_15 ^ t_15
lix_xor
  #(.W (32))
  u181_lix_xor
   (.i_x (u_15),
    .i_y (t_15),
    .o_z (z_15));



// u_16 ^ t_16
lix_xor
  #(.W (32))
  u182_lix_xor
   (.i_x (u_16),
    .i_y (t_16),
    .o_z (z_16));



// u_17 ^ t_17
lix_xor
  #(.W (32))
  u183_lix_xor
   (.i_x (u_17),
    .i_y (t_17),
    .o_z (z_17));



// u_18 ^ t_18
lix_xor
  #(.W (32))
  u184_lix_xor
   (.i_x (u_18),
    .i_y (t_18),
    .o_z (z_18));



// u_19 ^ t_19
lix_xor
  #(.W (32))
  u185_lix_xor
   (.i_x (u_19),
    .i_y (t_19),
    .o_z (z_19));



// z_1 ^ z_0
lix_xor
  #(.W (32))
  u186_lix_xor
   (.i_x (z_0),
    .i_y (z_1),
    .o_z (zxz_0));



// z_2 ^ zxz_0
lix_xor
  #(.W (32))
  u187_lix_xor
   (.i_x (z_2),
    .i_y (zxz_0),
    .o_z (zxz_1));



// z_3 ^ zxz_1
lix_xor
  #(.W (32))
  u188_lix_xor
   (.i_x (z_3),
    .i_y (zxz_1),
    .o_z (zxz_2));



// z_5 ^ z_4
lix_xor
  #(.W (32))
  u189_lix_xor
   (.i_x (z_4),
    .i_y (z_5),
    .o_z (zxz_3));



// z_6 ^ zxz_3
lix_xor
  #(.W (32))
  u190_lix_xor
   (.i_x (z_6),
    .i_y (zxz_3),
    .o_z (zxz_4));



// z_7 ^ zxz_4
lix_xor
  #(.W (32))
  u191_lix_xor
   (.i_x (z_7),
    .i_y (zxz_4),
    .o_z (zxz_5));



// z_9 ^ z_8
lix_xor
  #(.W (32))
  u192_lix_xor
   (.i_x (z_8),
    .i_y (z_9),
    .o_z (zxz_6));



// z_10 ^ zxz_6
lix_xor
  #(.W (32))
  u193_lix_xor
   (.i_x (z_10),
    .i_y (zxz_6),
    .o_z (zxz_7));



// z_11 ^ zxz_7
lix_xor
  #(.W (32))
  u194_lix_xor
   (.i_x (z_11),
    .i_y (zxz_7),
    .o_z (zxz_8));



// z_13 ^ z_12
lix_xor
  #(.W (32))
  u195_lix_xor
   (.i_x (z_12),
    .i_y (z_13),
    .o_z (zxz_9));



// z_14 ^ zxz_9
lix_xor
  #(.W (32))
  u196_lix_xor
   (.i_x (z_14),
    .i_y (zxz_9),
    .o_z (zxz_10));



// z_15 ^ zxz_10
lix_xor
  #(.W (32))
  u197_lix_xor
   (.i_x (z_15),
    .i_y (zxz_10),
    .o_z (zxz_11));



// z_17 ^ z_16
lix_xor
  #(.W (32))
  u198_lix_xor
   (.i_x (z_16),
    .i_y (z_17),
    .o_z (zxz_12));



// z_18 ^ zxz_12
lix_xor
  #(.W (32))
  u199_lix_xor
   (.i_x (z_18),
    .i_y (zxz_12),
    .o_z (zxz_13));



// z_19 ^ zxz_13
lix_xor
  #(.W (32))
  u200_lix_xor
   (.i_x (z_19),
    .i_y (zxz_13),
    .o_z (zxz_14));



// k_0 ^ zxz_2
lix_xor
  #(.W (32))
  u201_lix_xor
   (.i_x (k_0),
    .i_y (zxz_2),
    .o_z (o_c[0+:32]));



// k_1 ^ zxz_5
lix_xor
  #(.W (32))
  u202_lix_xor
   (.i_x (k_1),
    .i_y (zxz_5),
    .o_z (o_c[32+:32]));



// k_2 ^ zxz_8
lix_xor
  #(.W (32))
  u203_lix_xor
   (.i_x (k_2),
    .i_y (zxz_8),
    .o_z (o_c[64+:32]));



// k_3 ^ zxz_11
lix_xor
  #(.W (32))
  u204_lix_xor
   (.i_x (k_3),
    .i_y (zxz_11),
    .o_z (o_c[96+:32]));



// k_4 ^ zxz_14
lix_xor
  #(.W (32))
  u205_lix_xor
   (.i_x (k_4),
    .i_y (zxz_14),
    .o_z (o_c[128+:32]));



endmodule
