//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2024-04-26
// File Name     : ConvertAB_n2k32_0.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module ConvertAB_n2k32_0(
    input  wire         clk_i,
    input  wire         rst_ni,
    input  wire         i_dvld,
    input  wire         i_rvld,
    input  wire [319:0] i_n,
    input  wire  [63:0] i_a,
    output wire  [63:0] o_z);

wire     [31:0] x;
wire     [31:0] xd;
wire     [63:0] xp;
wire     [31:0] y;
wire     [31:0] yd;
wire     [63:0] yp;
wire            vrl;
wire            vy;

// ------------------------------------------------------------------------------
// Connect input port to left leaf data
// ------------------------------------------------------------------------------
assign x[ 0+:32] = i_a[ 0+:32];


// ------------------------------------------------------------------------------
// Connect left leaf data to Expand'input
// ------------------------------------------------------------------------------
assign xd[ 0+:32] = x[ 0+:32];


// ------------------------------------------------------------------------------
// Do a Expand(left leaf) instance
// ------------------------------------------------------------------------------
Expand1_n1o2k32
  u0_Expand1_n1o2k32
   (.i_x  (xd[0+:32]),
    .o_xp (xp[0+:64]));



// ------------------------------------------------------------------------------
// Connect i_dvld to right leaf valid
// ------------------------------------------------------------------------------
assign vrl = i_dvld;


// ------------------------------------------------------------------------------
// Connect input port to rifht leaf data
// ------------------------------------------------------------------------------
assign y[ 0+:32] = i_a[32+:32];


// ------------------------------------------------------------------------------
// Connect right leaf valid to right leaf output
// ------------------------------------------------------------------------------
assign vy = vrl;


// ------------------------------------------------------------------------------
// Connect right leaf data to Expand'input
// ------------------------------------------------------------------------------
assign yd[ 0+:32] = y[ 0+:32];


// ------------------------------------------------------------------------------
// Do a Expand(right leaf) instance
// ------------------------------------------------------------------------------
Expand2_n1o2k32
  u1_Expand2_n1o2k32
   (.i_x  (yd[0+:32]),
    .o_xp (yp[0+:64]));



// ------------------------------------------------------------------------------
// Do a KSA instance
// ------------------------------------------------------------------------------
SecKSA_n2k32_0
  u2_SecKSA_n2k32_0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (vy),
    .i_rvld (i_rvld),
    .i_n    (i_n[0+:320]),
    .i_x    (xp[0+:64]),
    .i_y    (yp[0+:64]),
    .o_z    (o_z[0+:64]));


endmodule
