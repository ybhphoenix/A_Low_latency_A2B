//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2024-04-26
// File Name     : ConvertAB_RCA_tb_n4k32.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module ConvertAB_RCA_tb_n4k32;

logic           clk_i;
logic           rst_ni;
logic           i_dvld;
logic           i_rvld;
logic   [247:0] i_n;
logic   [127:0] i_a;
logic   [127:0] o_z;
logic           o_dvld;
logic   [127:0] a;
logic           dvld;
logic    [31:0] A;
logic    [31:0] B;
logic    [31:0] A_d;
logic           pass;
logic           rvld;

initial
begin
  clk_i = 1'd0;
  forever #(10/2) clk_i = ~clk_i;
end


initial
begin
 rst_ni = 1'd0;
 #100;
 rst_ni = 1'd1;
end


initial
begin
  i_n = 248'd0;
  repeat (15) @(posedge clk_i);
  forever begin
    @(posedge clk_i);
    for(int i = 0 ; i < 248 ; i++)begin
      i_n[i] = $random;
    end
  end
end


initial
begin
  a = 128'd0;
  repeat (15) @(posedge clk_i);
  forever begin
    @(posedge clk_i);
    for(int i = 0 ; i < 4 ; i++)begin
      a[i*32+:32] = $random;
    end
  end
end


initial
begin
  dvld = 1'd0;
  repeat (16) @(posedge clk_i);
    dvld = 1'd1;
  repeat (500) @(posedge clk_i);
    dvld = 1'd0;
end


initial
begin
  rvld = 1'd0;
  repeat (16) @(posedge clk_i);
    rvld = 1'd1;
  repeat (624) @(posedge clk_i);
    rvld = 1'd0;
end

assign i_a[0+:32] = a[0+:32] - a[32+:32] - a[64+:32] - a[96+:32] ;
assign i_a[32+:32] = a[32+:32];
assign i_a[64+:32] = a[64+:32];
assign i_a[96+:32] = a[96+:32];
assign i_dvld = dvld;
assign i_rvld = rvld;
ConvertAB_RCA_n4k32_1
  dut_ConvertAB_RCA_n4k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n),
    .i_a    (i_a),
    .o_z    (o_z),
    .o_dvld (o_dvld));



assign A[0+:32] = i_a[0+:32] + i_a[32+:32] + i_a[64+:32] + i_a[96+:32] ;

assign B[0+:32] = o_z[0+:32] ^ o_z[32+:32] ^ o_z[64+:32] ^ o_z[96+:32] ;

reg  [31:0] shd_A_d [123:0];
always@(negedge rst_ni or posedge clk_i) begin
  if (~rst_ni)begin
    shd_A_d[0] <= 32'd0;
    shd_A_d[1] <= 32'd0;
    shd_A_d[2] <= 32'd0;
    shd_A_d[3] <= 32'd0;
    shd_A_d[4] <= 32'd0;
    shd_A_d[5] <= 32'd0;
    shd_A_d[6] <= 32'd0;
    shd_A_d[7] <= 32'd0;
    shd_A_d[8] <= 32'd0;
    shd_A_d[9] <= 32'd0;
    shd_A_d[10] <= 32'd0;
    shd_A_d[11] <= 32'd0;
    shd_A_d[12] <= 32'd0;
    shd_A_d[13] <= 32'd0;
    shd_A_d[14] <= 32'd0;
    shd_A_d[15] <= 32'd0;
    shd_A_d[16] <= 32'd0;
    shd_A_d[17] <= 32'd0;
    shd_A_d[18] <= 32'd0;
    shd_A_d[19] <= 32'd0;
    shd_A_d[20] <= 32'd0;
    shd_A_d[21] <= 32'd0;
    shd_A_d[22] <= 32'd0;
    shd_A_d[23] <= 32'd0;
    shd_A_d[24] <= 32'd0;
    shd_A_d[25] <= 32'd0;
    shd_A_d[26] <= 32'd0;
    shd_A_d[27] <= 32'd0;
    shd_A_d[28] <= 32'd0;
    shd_A_d[29] <= 32'd0;
    shd_A_d[30] <= 32'd0;
    shd_A_d[31] <= 32'd0;
    shd_A_d[32] <= 32'd0;
    shd_A_d[33] <= 32'd0;
    shd_A_d[34] <= 32'd0;
    shd_A_d[35] <= 32'd0;
    shd_A_d[36] <= 32'd0;
    shd_A_d[37] <= 32'd0;
    shd_A_d[38] <= 32'd0;
    shd_A_d[39] <= 32'd0;
    shd_A_d[40] <= 32'd0;
    shd_A_d[41] <= 32'd0;
    shd_A_d[42] <= 32'd0;
    shd_A_d[43] <= 32'd0;
    shd_A_d[44] <= 32'd0;
    shd_A_d[45] <= 32'd0;
    shd_A_d[46] <= 32'd0;
    shd_A_d[47] <= 32'd0;
    shd_A_d[48] <= 32'd0;
    shd_A_d[49] <= 32'd0;
    shd_A_d[50] <= 32'd0;
    shd_A_d[51] <= 32'd0;
    shd_A_d[52] <= 32'd0;
    shd_A_d[53] <= 32'd0;
    shd_A_d[54] <= 32'd0;
    shd_A_d[55] <= 32'd0;
    shd_A_d[56] <= 32'd0;
    shd_A_d[57] <= 32'd0;
    shd_A_d[58] <= 32'd0;
    shd_A_d[59] <= 32'd0;
    shd_A_d[60] <= 32'd0;
    shd_A_d[61] <= 32'd0;
    shd_A_d[62] <= 32'd0;
    shd_A_d[63] <= 32'd0;
    shd_A_d[64] <= 32'd0;
    shd_A_d[65] <= 32'd0;
    shd_A_d[66] <= 32'd0;
    shd_A_d[67] <= 32'd0;
    shd_A_d[68] <= 32'd0;
    shd_A_d[69] <= 32'd0;
    shd_A_d[70] <= 32'd0;
    shd_A_d[71] <= 32'd0;
    shd_A_d[72] <= 32'd0;
    shd_A_d[73] <= 32'd0;
    shd_A_d[74] <= 32'd0;
    shd_A_d[75] <= 32'd0;
    shd_A_d[76] <= 32'd0;
    shd_A_d[77] <= 32'd0;
    shd_A_d[78] <= 32'd0;
    shd_A_d[79] <= 32'd0;
    shd_A_d[80] <= 32'd0;
    shd_A_d[81] <= 32'd0;
    shd_A_d[82] <= 32'd0;
    shd_A_d[83] <= 32'd0;
    shd_A_d[84] <= 32'd0;
    shd_A_d[85] <= 32'd0;
    shd_A_d[86] <= 32'd0;
    shd_A_d[87] <= 32'd0;
    shd_A_d[88] <= 32'd0;
    shd_A_d[89] <= 32'd0;
    shd_A_d[90] <= 32'd0;
    shd_A_d[91] <= 32'd0;
    shd_A_d[92] <= 32'd0;
    shd_A_d[93] <= 32'd0;
    shd_A_d[94] <= 32'd0;
    shd_A_d[95] <= 32'd0;
    shd_A_d[96] <= 32'd0;
    shd_A_d[97] <= 32'd0;
    shd_A_d[98] <= 32'd0;
    shd_A_d[99] <= 32'd0;
    shd_A_d[100] <= 32'd0;
    shd_A_d[101] <= 32'd0;
    shd_A_d[102] <= 32'd0;
    shd_A_d[103] <= 32'd0;
    shd_A_d[104] <= 32'd0;
    shd_A_d[105] <= 32'd0;
    shd_A_d[106] <= 32'd0;
    shd_A_d[107] <= 32'd0;
    shd_A_d[108] <= 32'd0;
    shd_A_d[109] <= 32'd0;
    shd_A_d[110] <= 32'd0;
    shd_A_d[111] <= 32'd0;
    shd_A_d[112] <= 32'd0;
    shd_A_d[113] <= 32'd0;
    shd_A_d[114] <= 32'd0;
    shd_A_d[115] <= 32'd0;
    shd_A_d[116] <= 32'd0;
    shd_A_d[117] <= 32'd0;
    shd_A_d[118] <= 32'd0;
    shd_A_d[119] <= 32'd0;
    shd_A_d[120] <= 32'd0;
    shd_A_d[121] <= 32'd0;
    shd_A_d[122] <= 32'd0;
    shd_A_d[123] <= 32'd0;
  end else begin
    shd_A_d[0] <= A[0+:32];
    shd_A_d[1] <= shd_A_d[0];
    shd_A_d[2] <= shd_A_d[1];
    shd_A_d[3] <= shd_A_d[2];
    shd_A_d[4] <= shd_A_d[3];
    shd_A_d[5] <= shd_A_d[4];
    shd_A_d[6] <= shd_A_d[5];
    shd_A_d[7] <= shd_A_d[6];
    shd_A_d[8] <= shd_A_d[7];
    shd_A_d[9] <= shd_A_d[8];
    shd_A_d[10] <= shd_A_d[9];
    shd_A_d[11] <= shd_A_d[10];
    shd_A_d[12] <= shd_A_d[11];
    shd_A_d[13] <= shd_A_d[12];
    shd_A_d[14] <= shd_A_d[13];
    shd_A_d[15] <= shd_A_d[14];
    shd_A_d[16] <= shd_A_d[15];
    shd_A_d[17] <= shd_A_d[16];
    shd_A_d[18] <= shd_A_d[17];
    shd_A_d[19] <= shd_A_d[18];
    shd_A_d[20] <= shd_A_d[19];
    shd_A_d[21] <= shd_A_d[20];
    shd_A_d[22] <= shd_A_d[21];
    shd_A_d[23] <= shd_A_d[22];
    shd_A_d[24] <= shd_A_d[23];
    shd_A_d[25] <= shd_A_d[24];
    shd_A_d[26] <= shd_A_d[25];
    shd_A_d[27] <= shd_A_d[26];
    shd_A_d[28] <= shd_A_d[27];
    shd_A_d[29] <= shd_A_d[28];
    shd_A_d[30] <= shd_A_d[29];
    shd_A_d[31] <= shd_A_d[30];
    shd_A_d[32] <= shd_A_d[31];
    shd_A_d[33] <= shd_A_d[32];
    shd_A_d[34] <= shd_A_d[33];
    shd_A_d[35] <= shd_A_d[34];
    shd_A_d[36] <= shd_A_d[35];
    shd_A_d[37] <= shd_A_d[36];
    shd_A_d[38] <= shd_A_d[37];
    shd_A_d[39] <= shd_A_d[38];
    shd_A_d[40] <= shd_A_d[39];
    shd_A_d[41] <= shd_A_d[40];
    shd_A_d[42] <= shd_A_d[41];
    shd_A_d[43] <= shd_A_d[42];
    shd_A_d[44] <= shd_A_d[43];
    shd_A_d[45] <= shd_A_d[44];
    shd_A_d[46] <= shd_A_d[45];
    shd_A_d[47] <= shd_A_d[46];
    shd_A_d[48] <= shd_A_d[47];
    shd_A_d[49] <= shd_A_d[48];
    shd_A_d[50] <= shd_A_d[49];
    shd_A_d[51] <= shd_A_d[50];
    shd_A_d[52] <= shd_A_d[51];
    shd_A_d[53] <= shd_A_d[52];
    shd_A_d[54] <= shd_A_d[53];
    shd_A_d[55] <= shd_A_d[54];
    shd_A_d[56] <= shd_A_d[55];
    shd_A_d[57] <= shd_A_d[56];
    shd_A_d[58] <= shd_A_d[57];
    shd_A_d[59] <= shd_A_d[58];
    shd_A_d[60] <= shd_A_d[59];
    shd_A_d[61] <= shd_A_d[60];
    shd_A_d[62] <= shd_A_d[61];
    shd_A_d[63] <= shd_A_d[62];
    shd_A_d[64] <= shd_A_d[63];
    shd_A_d[65] <= shd_A_d[64];
    shd_A_d[66] <= shd_A_d[65];
    shd_A_d[67] <= shd_A_d[66];
    shd_A_d[68] <= shd_A_d[67];
    shd_A_d[69] <= shd_A_d[68];
    shd_A_d[70] <= shd_A_d[69];
    shd_A_d[71] <= shd_A_d[70];
    shd_A_d[72] <= shd_A_d[71];
    shd_A_d[73] <= shd_A_d[72];
    shd_A_d[74] <= shd_A_d[73];
    shd_A_d[75] <= shd_A_d[74];
    shd_A_d[76] <= shd_A_d[75];
    shd_A_d[77] <= shd_A_d[76];
    shd_A_d[78] <= shd_A_d[77];
    shd_A_d[79] <= shd_A_d[78];
    shd_A_d[80] <= shd_A_d[79];
    shd_A_d[81] <= shd_A_d[80];
    shd_A_d[82] <= shd_A_d[81];
    shd_A_d[83] <= shd_A_d[82];
    shd_A_d[84] <= shd_A_d[83];
    shd_A_d[85] <= shd_A_d[84];
    shd_A_d[86] <= shd_A_d[85];
    shd_A_d[87] <= shd_A_d[86];
    shd_A_d[88] <= shd_A_d[87];
    shd_A_d[89] <= shd_A_d[88];
    shd_A_d[90] <= shd_A_d[89];
    shd_A_d[91] <= shd_A_d[90];
    shd_A_d[92] <= shd_A_d[91];
    shd_A_d[93] <= shd_A_d[92];
    shd_A_d[94] <= shd_A_d[93];
    shd_A_d[95] <= shd_A_d[94];
    shd_A_d[96] <= shd_A_d[95];
    shd_A_d[97] <= shd_A_d[96];
    shd_A_d[98] <= shd_A_d[97];
    shd_A_d[99] <= shd_A_d[98];
    shd_A_d[100] <= shd_A_d[99];
    shd_A_d[101] <= shd_A_d[100];
    shd_A_d[102] <= shd_A_d[101];
    shd_A_d[103] <= shd_A_d[102];
    shd_A_d[104] <= shd_A_d[103];
    shd_A_d[105] <= shd_A_d[104];
    shd_A_d[106] <= shd_A_d[105];
    shd_A_d[107] <= shd_A_d[106];
    shd_A_d[108] <= shd_A_d[107];
    shd_A_d[109] <= shd_A_d[108];
    shd_A_d[110] <= shd_A_d[109];
    shd_A_d[111] <= shd_A_d[110];
    shd_A_d[112] <= shd_A_d[111];
    shd_A_d[113] <= shd_A_d[112];
    shd_A_d[114] <= shd_A_d[113];
    shd_A_d[115] <= shd_A_d[114];
    shd_A_d[116] <= shd_A_d[115];
    shd_A_d[117] <= shd_A_d[116];
    shd_A_d[118] <= shd_A_d[117];
    shd_A_d[119] <= shd_A_d[118];
    shd_A_d[120] <= shd_A_d[119];
    shd_A_d[121] <= shd_A_d[120];
    shd_A_d[122] <= shd_A_d[121];
    shd_A_d[123] <= shd_A_d[122];
  end
end
assign A_d[31:0] = shd_A_d[123];


assign pass = B[ 0+:32]  ==  A_d[ 0+:32];


logic fail;
initial
begin
  fail = 1'd0;
  forever begin
    @(posedge clk_i);
    if (pass != 1'd1 && o_dvld == 1'd1)begin
       $display("Test_Failed");
       fail = 1'd1;
    end
  end
end

initial
begin
  #7000;
  @(posedge clk_i);
  if (fail == 1'b0)begin
    $display("Test_Passed");
  end
end


initial
begin
  #8000;
  $finish;
end

endmodule
