//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2023-10-08
// File Name     : SecAnd_PINI1_n3k1_1.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecAnd_PINI1_n3k1_1(
    input  wire       clk_i,
    input  wire       rst_ni,
    input  wire       i_dvld,
    input  wire       i_rvld,
    input  wire [2:0] i_n,
    input  wire [2:0] i_x,
    input  wire [2:0] i_y,
    output wire [2:0] o_c,
    output wire       o_dvld);

(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire  vldd1;// synopsys keep_signal_name "vldd1" 
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xd_0;// synopsys keep_signal_name "xd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xd_1;// synopsys keep_signal_name "xd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xd_2;// synopsys keep_signal_name "xd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yd_0;// synopsys keep_signal_name "yd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yd_1;// synopsys keep_signal_name "yd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yd_2;// synopsys keep_signal_name "yd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_0;// synopsys keep_signal_name "r_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_1;// synopsys keep_signal_name "r_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_2;// synopsys keep_signal_name "r_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_3;// synopsys keep_signal_name "r_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_4;// synopsys keep_signal_name "r_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] r_5;// synopsys keep_signal_name "r_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_0;// synopsys keep_signal_name "yxn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_1;// synopsys keep_signal_name "yxn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_2;// synopsys keep_signal_name "yxn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_3;// synopsys keep_signal_name "yxn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_4;// synopsys keep_signal_name "yxn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] yxn_5;// synopsys keep_signal_name "yxn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_0;// synopsys keep_signal_name "v_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_1;// synopsys keep_signal_name "v_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_2;// synopsys keep_signal_name "v_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_3;// synopsys keep_signal_name "v_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_4;// synopsys keep_signal_name "v_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] v_5;// synopsys keep_signal_name "v_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire vldd2;
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_0;// synopsys keep_signal_name "xdn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_1;// synopsys keep_signal_name "xdn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_2;// synopsys keep_signal_name "xdn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_3;// synopsys keep_signal_name "xdn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_4;// synopsys keep_signal_name "xdn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xdn_5;// synopsys keep_signal_name "xdn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_0;// synopsys keep_signal_name "xar_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_1;// synopsys keep_signal_name "xar_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_2;// synopsys keep_signal_name "xar_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_3;// synopsys keep_signal_name "xar_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_4;// synopsys keep_signal_name "xar_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xar_5;// synopsys keep_signal_name "xar_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_0;// synopsys keep_signal_name "u_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_1;// synopsys keep_signal_name "u_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_2;// synopsys keep_signal_name "u_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_3;// synopsys keep_signal_name "u_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_4;// synopsys keep_signal_name "u_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] u_5;// synopsys keep_signal_name "u_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xay_0;// synopsys keep_signal_name "xay_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xay_1;// synopsys keep_signal_name "xay_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xay_2;// synopsys keep_signal_name "xay_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] k_0;// synopsys keep_signal_name "k_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] k_1;// synopsys keep_signal_name "k_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] k_2;// synopsys keep_signal_name "k_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_0;// synopsys keep_signal_name "xav_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_1;// synopsys keep_signal_name "xav_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_2;// synopsys keep_signal_name "xav_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_3;// synopsys keep_signal_name "xav_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_4;// synopsys keep_signal_name "xav_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] xav_5;// synopsys keep_signal_name "xav_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_0;// synopsys keep_signal_name "t_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_1;// synopsys keep_signal_name "t_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_2;// synopsys keep_signal_name "t_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_3;// synopsys keep_signal_name "t_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_4;// synopsys keep_signal_name "t_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] t_5;// synopsys keep_signal_name "t_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_0;// synopsys keep_signal_name "z_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_1;// synopsys keep_signal_name "z_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_2;// synopsys keep_signal_name "z_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_3;// synopsys keep_signal_name "z_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_4;// synopsys keep_signal_name "z_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] z_5;// synopsys keep_signal_name "z_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] zxz_0;// synopsys keep_signal_name "zxz_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] zxz_1;// synopsys keep_signal_name "zxz_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [0:0] zxz_2;// synopsys keep_signal_name "zxz_2"

// delay i_dvld
lix_reg
  #(.W (1))
  u0_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (i_dvld),
    .o_z    (vldd1));



// delay i_x[0+:1]
lix_reg
  #(.W (1))
  u1_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[0+:1]),
    .o_z    (xd_0));



// delay i_x[1+:1]
lix_reg
  #(.W (1))
  u2_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[1+:1]),
    .o_z    (xd_1));



// delay i_x[2+:1]
lix_reg
  #(.W (1))
  u3_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[2+:1]),
    .o_z    (xd_2));



// delay i_y[0+:1]
lix_reg
  #(.W (1))
  u4_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[0+:1]),
    .o_z    (yd_0));



// delay i_y[1+:1]
lix_reg
  #(.W (1))
  u5_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[1+:1]),
    .o_z    (yd_1));



// delay i_y[2+:1]
lix_reg
  #(.W (1))
  u6_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[2+:1]),
    .o_z    (yd_2));



// delay i_n0
lix_reg
  #(.W (1))
  u7_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:1]),
    .o_z    (r_0));



// delay i_n1
lix_reg
  #(.W (1))
  u8_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[1+:1]),
    .o_z    (r_1));



// delay i_n0
lix_reg
  #(.W (1))
  u9_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:1]),
    .o_z    (r_2));



// delay i_n2
lix_reg
  #(.W (1))
  u10_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[2+:1]),
    .o_z    (r_3));



// delay i_n1
lix_reg
  #(.W (1))
  u11_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[1+:1]),
    .o_z    (r_4));



// delay i_n2
lix_reg
  #(.W (1))
  u12_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[2+:1]),
    .o_z    (r_5));



// i_y[0+:1] ^ i_n[0+:1]
lix_xor
  #(.W (1))
  u13_lix_xor
   (.i_x (i_y[1+:1]),
    .i_y (i_n[0+:1]),
    .o_z (yxn_0));



// i_y[0+:1] ^ i_n[1+:1]
lix_xor
  #(.W (1))
  u14_lix_xor
   (.i_x (i_y[2+:1]),
    .i_y (i_n[1+:1]),
    .o_z (yxn_1));



// i_y[1+:1] ^ i_n[0+:1]
lix_xor
  #(.W (1))
  u15_lix_xor
   (.i_x (i_y[0+:1]),
    .i_y (i_n[0+:1]),
    .o_z (yxn_2));



// i_y[1+:1] ^ i_n[2+:1]
lix_xor
  #(.W (1))
  u16_lix_xor
   (.i_x (i_y[2+:1]),
    .i_y (i_n[2+:1]),
    .o_z (yxn_3));



// i_y[2+:1] ^ i_n[1+:1]
lix_xor
  #(.W (1))
  u17_lix_xor
   (.i_x (i_y[0+:1]),
    .i_y (i_n[1+:1]),
    .o_z (yxn_4));



// i_y[2+:1] ^ i_n[2+:1]
lix_xor
  #(.W (1))
  u18_lix_xor
   (.i_x (i_y[1+:1]),
    .i_y (i_n[2+:1]),
    .o_z (yxn_5));



// delay yxn_0
lix_reg
  #(.W (1))
  u19_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_0),
    .o_z    (v_0));



// delay yxn_1
lix_reg
  #(.W (1))
  u20_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_1),
    .o_z    (v_1));



// delay yxn_2
lix_reg
  #(.W (1))
  u21_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_2),
    .o_z    (v_2));



// delay yxn_3
lix_reg
  #(.W (1))
  u22_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_3),
    .o_z    (v_3));



// delay yxn_4
lix_reg
  #(.W (1))
  u23_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_4),
    .o_z    (v_4));



// delay yxn_5
lix_reg
  #(.W (1))
  u24_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_5),
    .o_z    (v_5));



// delay vldd1
lix_reg
  #(.W (1))
  u25_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (vldd1),
    .o_z    (vldd2));



// not  xd_0
lix_not
  #(.W (1))
  u26_lix_not
   (.i_x (xd_0),
    .o_z (xdn_0));



// not  xd_1
lix_not
  #(.W (1))
  u27_lix_not
   (.i_x (xd_1),
    .o_z (xdn_1));



// not  xd_2
lix_not
  #(.W (1))
  u28_lix_not
   (.i_x (xd_2),
    .o_z (xdn_2));



// ~xd_0 & r_0
lix_and
  #(.W (1))
  u29_lix_and
   (.i_x (xdn_0),
    .i_y (r_0),
    .o_z (xar_0));



// ~xd_0 & r_1
lix_and
  #(.W (1))
  u30_lix_and
   (.i_x (xdn_0),
    .i_y (r_1),
    .o_z (xar_1));



// ~xd_1 & r_2
lix_and
  #(.W (1))
  u31_lix_and
   (.i_x (xdn_1),
    .i_y (r_2),
    .o_z (xar_2));



// ~xd_1 & r_3
lix_and
  #(.W (1))
  u32_lix_and
   (.i_x (xdn_1),
    .i_y (r_3),
    .o_z (xar_3));



// ~xd_2 & r_4
lix_and
  #(.W (1))
  u33_lix_and
   (.i_x (xdn_2),
    .i_y (r_4),
    .o_z (xar_4));



// ~xd_2 & r_5
lix_and
  #(.W (1))
  u34_lix_and
   (.i_x (xdn_2),
    .i_y (r_5),
    .o_z (xar_5));



// delay ~xd_0 & r_0
lix_reg
  #(.W (1))
  u35_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_0),
    .o_z    (u_0));



// delay ~xd_1 & r_1
lix_reg
  #(.W (1))
  u36_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_1),
    .o_z    (u_1));



// delay ~xd_2 & r_2
lix_reg
  #(.W (1))
  u37_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_2),
    .o_z    (u_2));



// delay ~xd_3 & r_3
lix_reg
  #(.W (1))
  u38_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_3),
    .o_z    (u_3));



// delay ~xd_4 & r_4
lix_reg
  #(.W (1))
  u39_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_4),
    .o_z    (u_4));



// delay ~xd_5 & r_5
lix_reg
  #(.W (1))
  u40_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_5),
    .o_z    (u_5));



// xd_0 & yd_0
lix_and
  #(.W (1))
  u41_lix_and
   (.i_x (xd_0),
    .i_y (yd_0),
    .o_z (xay_0));



// xd_1 & yd_1
lix_and
  #(.W (1))
  u42_lix_and
   (.i_x (xd_1),
    .i_y (yd_1),
    .o_z (xay_1));



// xd_2 & yd_2
lix_and
  #(.W (1))
  u43_lix_and
   (.i_x (xd_2),
    .i_y (yd_2),
    .o_z (xay_2));



// delay xd_0 & yd_0
lix_reg
  #(.W (1))
  u44_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_0),
    .o_z    (k_0));



// delay xd_1 & yd_1
lix_reg
  #(.W (1))
  u45_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_1),
    .o_z    (k_1));



// delay xd_2 & yd_2
lix_reg
  #(.W (1))
  u46_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_2),
    .o_z    (k_2));



// xd_0 & v_0
lix_and
  #(.W (1))
  u47_lix_and
   (.i_x (xd_0),
    .i_y (v_0),
    .o_z (xav_0));



// xd_0 & v_1
lix_and
  #(.W (1))
  u48_lix_and
   (.i_x (xd_0),
    .i_y (v_1),
    .o_z (xav_1));



// xd_1 & v_2
lix_and
  #(.W (1))
  u49_lix_and
   (.i_x (xd_1),
    .i_y (v_2),
    .o_z (xav_2));



// xd_1 & v_3
lix_and
  #(.W (1))
  u50_lix_and
   (.i_x (xd_1),
    .i_y (v_3),
    .o_z (xav_3));



// xd_2 & v_4
lix_and
  #(.W (1))
  u51_lix_and
   (.i_x (xd_2),
    .i_y (v_4),
    .o_z (xav_4));



// xd_2 & v_5
lix_and
  #(.W (1))
  u52_lix_and
   (.i_x (xd_2),
    .i_y (v_5),
    .o_z (xav_5));



// delay xd_0 & v_0
lix_reg
  #(.W (1))
  u53_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_0),
    .o_z    (t_0));



// delay xd_1 & v_1
lix_reg
  #(.W (1))
  u54_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_1),
    .o_z    (t_1));



// delay xd_2 & v_2
lix_reg
  #(.W (1))
  u55_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_2),
    .o_z    (t_2));



// delay xd_3 & v_3
lix_reg
  #(.W (1))
  u56_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_3),
    .o_z    (t_3));



// delay xd_4 & v_4
lix_reg
  #(.W (1))
  u57_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_4),
    .o_z    (t_4));



// delay xd_5 & v_5
lix_reg
  #(.W (1))
  u58_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_5),
    .o_z    (t_5));



// u_0 ^ t_0
lix_xor
  #(.W (1))
  u59_lix_xor
   (.i_x (u_0),
    .i_y (t_0),
    .o_z (z_0));



// u_1 ^ t_1
lix_xor
  #(.W (1))
  u60_lix_xor
   (.i_x (u_1),
    .i_y (t_1),
    .o_z (z_1));



// u_2 ^ t_2
lix_xor
  #(.W (1))
  u61_lix_xor
   (.i_x (u_2),
    .i_y (t_2),
    .o_z (z_2));



// u_3 ^ t_3
lix_xor
  #(.W (1))
  u62_lix_xor
   (.i_x (u_3),
    .i_y (t_3),
    .o_z (z_3));



// u_4 ^ t_4
lix_xor
  #(.W (1))
  u63_lix_xor
   (.i_x (u_4),
    .i_y (t_4),
    .o_z (z_4));



// u_5 ^ t_5
lix_xor
  #(.W (1))
  u64_lix_xor
   (.i_x (u_5),
    .i_y (t_5),
    .o_z (z_5));



// z_1 ^ z_0
lix_xor
  #(.W (1))
  u65_lix_xor
   (.i_x (z_0),
    .i_y (z_1),
    .o_z (zxz_0));



// z_3 ^ z_2
lix_xor
  #(.W (1))
  u66_lix_xor
   (.i_x (z_2),
    .i_y (z_3),
    .o_z (zxz_1));



// z_5 ^ z_4
lix_xor
  #(.W (1))
  u67_lix_xor
   (.i_x (z_4),
    .i_y (z_5),
    .o_z (zxz_2));



// k_0 ^ zxz_0
lix_xor
  #(.W (1))
  u68_lix_xor
   (.i_x (k_0),
    .i_y (zxz_0),
    .o_z (o_c[0+:1]));



// k_1 ^ zxz_1
lix_xor
  #(.W (1))
  u69_lix_xor
   (.i_x (k_1),
    .i_y (zxz_1),
    .o_z (o_c[1+:1]));



// k_2 ^ zxz_2
lix_xor
  #(.W (1))
  u70_lix_xor
   (.i_x (k_2),
    .i_y (zxz_2),
    .o_z (o_c[2+:1]));



assign o_dvld = vldd2;

endmodule
