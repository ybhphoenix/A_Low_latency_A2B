//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2023-10-08
// File Name     : SecKSA_1l_n4k32.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecKSA_1l_n4k32   #(
    parameter  SHIFT = 1,
    parameter  POW = 2**SHIFT
  )(
    input  wire         clk_i,
    input  wire         rst_ni,
    input  wire         i_dvld,
    input  wire         i_rvld,
    input  wire [383:0] i_n,
    input  wire [127:0] i_p,
    input  wire [127:0] i_g,
    output wire [127:0] o_p,
    output wire [127:0] o_g,
    output wire         o_dvld);

wire    [127:0] tmp1;
wire    [127:0] a1;
wire    [127:0] gd;
wire    [127:0] tmp2;
wire    [127:0] a2;

// ------------------------------------------------------------------------------
// tmp[i]=(g[i]<<pow)&MASK;
// ------------------------------------------------------------------------------
assign tmp1[  0+: 32] = i_g[  0+: 32]  <<  POW;
assign tmp1[ 32+: 32] = i_g[ 32+: 32]  <<  POW;
assign tmp1[ 64+: 32] = i_g[ 64+: 32]  <<  POW;
assign tmp1[ 96+: 32] = i_g[ 96+: 32]  <<  POW;


// ------------------------------------------------------------------------------
// tmp[i]=(p[i]<<pow)&MASK;
// ------------------------------------------------------------------------------
assign tmp2[  0+: 32] = i_p[  0+: 32]  <<  POW;
assign tmp2[ 32+: 32] = i_p[ 32+: 32]  <<  POW;
assign tmp2[ 64+: 32] = i_p[ 64+: 32]  <<  POW;
assign tmp2[ 96+: 32] = i_p[ 96+: 32]  <<  POW;


// ------------------------------------------------------------------------------
// SecAnd_PINI1(p,tmp,a,k,n);
// ------------------------------------------------------------------------------
SecAnd_PINI1_n4k32_1
  u0_SecAnd_PINI1_n4k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[0+:192]),
    .i_x    (i_p),
    .i_y    (tmp1),
    .o_c    (a1),
    .o_dvld (o_dvld));



// ------------------------------------------------------------------------------
// SecAnd_PINI1(p,tmp,a,k,n);
// ------------------------------------------------------------------------------
SecAnd_PINI1_n4k32_0
  u1_SecAnd_PINI1_n4k32_0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[192+:192]),
    .i_x    (i_p),
    .i_y    (tmp2),
    .o_c    (a2));



// ------------------------------------------------------------------------------
// Delay i_g
// ------------------------------------------------------------------------------
lix_shr0
  #(.W (128),
    .N (2))
  u2_lix_shr0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_g),
    .o_z    (gd));



// ------------------------------------------------------------------------------
// g[i]=g[i]^a[i];
// ------------------------------------------------------------------------------
lix_xor
  #(.W (128))
  u3_lix_xor
   (.i_x (gd),
    .i_y (a1),
    .o_z (o_g));



// ------------------------------------------------------------------------------
// Connect a2 to output
// ------------------------------------------------------------------------------
assign o_p[  0+:128] = a2[  0+:128];

endmodule
