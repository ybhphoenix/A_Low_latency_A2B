//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2023-10-08
// File Name     : ConvertAB_n5k32_1.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module ConvertAB_n5k32_1(
    input  wire          clk_i,
    input  wire          rst_ni,
    input  wire          i_dvld,
    input  wire          i_rvld,
    input  wire [4799:0] i_n,
    input  wire  [159:0] i_a,
    output wire  [159:0] o_z,
    output wire          o_dvld);

wire     [63:0] x;
wire     [63:0] xd;
wire    [159:0] xp;
wire     [95:0] y;
wire     [95:0] yd;
wire    [159:0] yp;
wire            vrl;
wire            vy;
wire            vll;

// ------------------------------------------------------------------------------
// Do ConvertAB(left leaf) instance
// ------------------------------------------------------------------------------
ConvertAB_n2k32_1
  u0_ConvertAB_n2k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[0+:320]),
    .i_a    (i_a[0+:64]),
    .o_z    (x[0+:64]),
    .o_dvld (vll));



// ------------------------------------------------------------------------------
// Delay left leaf
// ------------------------------------------------------------------------------
lix_shr0
  #(.W (64),
    .N (12))
  u1_lix_shr0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vll),
    .i_en   (i_rvld),
    .i_x    (x[0+:64]),
    .o_z    (xd[0+:64]));



// ------------------------------------------------------------------------------
// Do a Expand(left leaf) instance
// ------------------------------------------------------------------------------
Expand1_n2o5k32
  u2_Expand1_n2o5k32
   (.i_x  (xd[0+:64]),
    .o_xp (xp[0+:160]));



// ------------------------------------------------------------------------------
// Do ConvertAB(right leaf) instance
// ------------------------------------------------------------------------------
ConvertAB_n3k32_1
  u3_ConvertAB_n3k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[320+:1280]),
    .i_a    (i_a[64+:96]),
    .o_z    (y[0+:96]),
    .o_dvld (vrl));



// ------------------------------------------------------------------------------
// Connect right leaf valid to right leaf output
// ------------------------------------------------------------------------------
assign vy = vrl;


// ------------------------------------------------------------------------------
// Connect right leaf data to Expand'input
// ------------------------------------------------------------------------------
assign yd[ 0+:96] = y[ 0+:96];


// ------------------------------------------------------------------------------
// Do a Expand(right leaf) instance
// ------------------------------------------------------------------------------
Expand2_n3o5k32
  u4_Expand2_n3o5k32
   (.i_x  (yd[0+:96]),
    .o_xp (yp[0+:160]));



// ------------------------------------------------------------------------------
// Do a KSA instance
// ------------------------------------------------------------------------------
SecKSA_n5k32_1
  u5_SecKSA_n5k32_1
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (vy),
    .i_rvld (i_rvld),
    .i_n    (i_n[1600+:3200]),
    .i_x    (xp[0+:160]),
    .i_y    (yp[0+:160]),
    .o_z    (o_z[0+:160]),
    .o_dvld (o_dvld));


endmodule
