//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2024-04-26
// File Name     : SecCSATree_n5k32.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecCSATree_n5k32(
    input  wire         clk_i,
    input  wire         rst_ni,
    input  wire         i_dvld,
    input  wire         i_rvld,
    input  wire [607:0] i_n,
    input  wire [159:0] i_x,
    output wire [159:0] o_s,
    output wire [159:0] o_c,
    output wire         o_dvld);

wire    [159:0] y1;
wire    [159:0] y2;
wire    [159:0] y3;
wire            vc;
wire     [31:0] xd;
wire    [127:0] s;
wire    [127:0] c;

// ------------------------------------------------------------------------------
// Do SecCSAtree instance
// ------------------------------------------------------------------------------
SecCSATree_n4k32
  u0_SecCSATree_n4k32
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (i_dvld),
    .i_rvld (i_rvld),
    .i_n    (i_n[0+:288]),
    .i_x    (i_x[0+:128]),
    .o_s    (s),
    .o_c    (c),
    .o_dvld (vc));



// ------------------------------------------------------------------------------
// Do pipeline instance
// ------------------------------------------------------------------------------
lix_shr0
  #(.W (32),
    .N (4))
  u1_lix_shr0
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[128+:32]),
    .o_z    (xd[0+:32]));



// ------------------------------------------------------------------------------
// for(i=0;i<n-1;i++) y1[i]=s[i];
// y1[n-1]=0;
// ------------------------------------------------------------------------------
assign y1[0+:32] = s[0+:32];
assign y1[32+:32] = s[32+:32];
assign y1[64+:32] = s[64+:32];
assign y1[96+:32] = s[96+:32];
assign y1[128+:32] = 32'd0;

// ------------------------------------------------------------------------------
// for(i=0;i<n-1;i++) y2[i]=c[i];
// y2[n-1]=0;
// ------------------------------------------------------------------------------
assign y2[0+:32] = c[0+:32];
assign y2[32+:32] = c[32+:32];
assign y2[64+:32] = c[64+:32];
assign y2[96+:32] = c[96+:32];
assign y2[128+:32] = 32'd0;

// ------------------------------------------------------------------------------
// for(i=0;i<n-1;i++) y3[i]=0;
// y3[n-1]=x[n-1];
// ------------------------------------------------------------------------------
assign y3[0+:32] = 32'd0;
assign y3[32+:32] = 32'd0;
assign y3[64+:32] = 32'd0;
assign y3[96+:32] = 32'd0;
assign y3[128+:32] = xd[0+:32];

// ------------------------------------------------------------------------------
// Do SecCSA instance
// ------------------------------------------------------------------------------
SecCSA_n5k32
  u2_SecCSA_n5k32
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_dvld (vc),
    .i_rvld (i_rvld),
    .i_n    (i_n[288+:320]),
    .i_x    (y1),
    .i_y    (y2),
    .i_c_in (y3),
    .o_s    (o_s),
    .o_c    (o_c),
    .o_dvld (o_dvld));


endmodule
